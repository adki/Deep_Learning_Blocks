
   dpu #(.P_DATA_TYPE    (DATA_TYPE )
        ,.P_DATA_WIDTH   (DATA_WIDTH)
        `ifdef DATA_FIXED_POINT
        ,.P_DATA_WIDTH_Q (DATA_WIDTH_Q)
        `endif
        ,.S_AXI_WIDTH_ID (P_AXI_WIDTH_SID)
        ,.S_AXI_WIDTH_AD (P_AXI_WIDTH_AD )
        ,.S_AXI_WIDTH_DA (P_AXI_WIDTH_DA )
        ,.M_AXI_WIDTH_ID (P_AXI_WIDTH_ID )
        ,.M_AXI_WIDTH_AD (P_AXI_WIDTH_AD )
        ,.M_AXI_WIDTH_DA (P_AXI_WIDTH_DA )
        ,.P_ADDR_BASE_CONF  (`DPU_ADDR_BASE_CONF  ),.P_SIZE_CONF  (`DPU_SIZE_CONF  )
        ,.P_ADDR_BASE_CONV  (`DPU_ADDR_BASE_CONV  ),.P_SIZE_CONV  (`DPU_SIZE_CONV  )
        ,.P_ADDR_BASE_POOL  (`DPU_ADDR_BASE_POOL  ),.P_SIZE_POOL  (`DPU_SIZE_POOL  )
        ,.P_ADDR_BASE_LINEAR(`DPU_ADDR_BASE_LINEAR),.P_SIZE_LINEAR(`DPU_SIZE_LINEAR)
        ,.P_ADDR_BASE_MOVER (`DPU_ADDR_BASE_MOVER ),.P_SIZE_MOVER (`DPU_SIZE_MOVER )
        ,.P_ADDR_BASE_DPU   (`DPU_ADDR_BASE_DPU   ),.P_SIZE_DPU   (`DPU_SIZE_DPU   ))
    u_dpu (
          .ARESETn                     ( ARESETn          )
        , .ACLK                        ( ACLK             )

        , .s_axi_AWID                  ( s_axi_AWID   [1] )
        , .s_axi_AWADDR                ( s_axi_AWADDR [1] )
        , .s_axi_AWLEN                 ( s_axi_AWLEN  [1] )
        , .s_axi_AWSIZE                ( s_axi_AWSIZE [1] )
        , .s_axi_AWBURST               ( s_axi_AWBURST[1] )
        , .s_axi_AWVALID               ( s_axi_AWVALID[1] )
        , .s_axi_AWREADY               ( s_axi_AWREADY[1] )
        , .s_axi_WDATA                 ( s_axi_WDATA  [1] )
        , .s_axi_WSTRB                 ( s_axi_WSTRB  [1] )
        , .s_axi_WLAST                 ( s_axi_WLAST  [1] )
        , .s_axi_WVALID                ( s_axi_WVALID [1] )
        , .s_axi_WREADY                ( s_axi_WREADY [1] )
        , .s_axi_BID                   ( s_axi_BID    [1] )
        , .s_axi_BRESP                 ( s_axi_BRESP  [1] )
        , .s_axi_BVALID                ( s_axi_BVALID [1] )
        , .s_axi_BREADY                ( s_axi_BREADY [1] )
        , .s_axi_ARID                  ( s_axi_ARID   [1] )
        , .s_axi_ARADDR                ( s_axi_ARADDR [1] )
        , .s_axi_ARLEN                 ( s_axi_ARLEN  [1] )
        , .s_axi_ARSIZE                ( s_axi_ARSIZE [1] )
        , .s_axi_ARBURST               ( s_axi_ARBURST[1] )
        , .s_axi_ARVALID               ( s_axi_ARVALID[1] )
        , .s_axi_ARREADY               ( s_axi_ARREADY[1] )
        , .s_axi_RID                   ( s_axi_RID    [1] )
        , .s_axi_RDATA                 ( s_axi_RDATA  [1] )
        , .s_axi_RRESP                 ( s_axi_RRESP  [1] )
        , .s_axi_RLAST                 ( s_axi_RLAST  [1] )
        , .s_axi_RVALID                ( s_axi_RVALID [1] )
        , .s_axi_RREADY                ( s_axi_RREADY [1] )

        , .m_axi_conv_rst_AWID         ( m_axi_AWID   [1] )
        , .m_axi_conv_rst_AWADDR       ( m_axi_AWADDR [1] )
        , .m_axi_conv_rst_AWLEN        ( m_axi_AWLEN  [1] )
        , .m_axi_conv_rst_AWSIZE       ( m_axi_AWSIZE [1] )
        , .m_axi_conv_rst_AWBURST      ( m_axi_AWBURST[1] )
        , .m_axi_conv_rst_AWVALID      ( m_axi_AWVALID[1] )
        , .m_axi_conv_rst_AWREADY      ( m_axi_AWREADY[1] )
        , .m_axi_conv_rst_WDATA        ( m_axi_WDATA  [1] )
        , .m_axi_conv_rst_WSTRB        ( m_axi_WSTRB  [1] )
        , .m_axi_conv_rst_WLAST        ( m_axi_WLAST  [1] )
        , .m_axi_conv_rst_WVALID       ( m_axi_WVALID [1] )
        , .m_axi_conv_rst_WREADY       ( m_axi_WREADY [1] )
        , .m_axi_conv_rst_BID          ( m_axi_BID    [1] )
        , .m_axi_conv_rst_BRESP        ( m_axi_BRESP  [1] )
        , .m_axi_conv_rst_BVALID       ( m_axi_BVALID [1] )
        , .m_axi_conv_rst_BREADY       ( m_axi_BREADY [1] )
        , .m_axi_conv_rst_ARID         ( m_axi_ARID   [1] )
        , .m_axi_conv_rst_ARADDR       ( m_axi_ARADDR [1] )
        , .m_axi_conv_rst_ARLEN        ( m_axi_ARLEN  [1] )
        , .m_axi_conv_rst_ARSIZE       ( m_axi_ARSIZE [1] )
        , .m_axi_conv_rst_ARBURST      ( m_axi_ARBURST[1] )
        , .m_axi_conv_rst_ARVALID      ( m_axi_ARVALID[1] )
        , .m_axi_conv_rst_ARREADY      ( m_axi_ARREADY[1] )
        , .m_axi_conv_rst_RID          ( m_axi_RID    [1] )
        , .m_axi_conv_rst_RDATA        ( m_axi_RDATA  [1] )
        , .m_axi_conv_rst_RRESP        ( m_axi_RRESP  [1] )
        , .m_axi_conv_rst_RLAST        ( m_axi_RLAST  [1] )
        , .m_axi_conv_rst_RVALID       ( m_axi_RVALID [1] )
        , .m_axi_conv_rst_RREADY       ( m_axi_RREADY [1] )

        , .m_axi_conv_knl_AWID         ( m_axi_AWID   [2] )
        , .m_axi_conv_knl_AWADDR       ( m_axi_AWADDR [2] )
        , .m_axi_conv_knl_AWLEN        ( m_axi_AWLEN  [2] )
        , .m_axi_conv_knl_AWSIZE       ( m_axi_AWSIZE [2] )
        , .m_axi_conv_knl_AWBURST      ( m_axi_AWBURST[2] )
        , .m_axi_conv_knl_AWVALID      ( m_axi_AWVALID[2] )
        , .m_axi_conv_knl_AWREADY      ( m_axi_AWREADY[2] )
        , .m_axi_conv_knl_WDATA        ( m_axi_WDATA  [2] )
        , .m_axi_conv_knl_WSTRB        ( m_axi_WSTRB  [2] )
        , .m_axi_conv_knl_WLAST        ( m_axi_WLAST  [2] )
        , .m_axi_conv_knl_WVALID       ( m_axi_WVALID [2] )
        , .m_axi_conv_knl_WREADY       ( m_axi_WREADY [2] )
        , .m_axi_conv_knl_BID          ( m_axi_BID    [2] )
        , .m_axi_conv_knl_BRESP        ( m_axi_BRESP  [2] )
        , .m_axi_conv_knl_BVALID       ( m_axi_BVALID [2] )
        , .m_axi_conv_knl_BREADY       ( m_axi_BREADY [2] )
        , .m_axi_conv_knl_ARID         ( m_axi_ARID   [2] )
        , .m_axi_conv_knl_ARADDR       ( m_axi_ARADDR [2] )
        , .m_axi_conv_knl_ARLEN        ( m_axi_ARLEN  [2] )
        , .m_axi_conv_knl_ARSIZE       ( m_axi_ARSIZE [2] )
        , .m_axi_conv_knl_ARBURST      ( m_axi_ARBURST[2] )
        , .m_axi_conv_knl_ARVALID      ( m_axi_ARVALID[2] )
        , .m_axi_conv_knl_ARREADY      ( m_axi_ARREADY[2] )
        , .m_axi_conv_knl_RID          ( m_axi_RID    [2] )
        , .m_axi_conv_knl_RDATA        ( m_axi_RDATA  [2] )
        , .m_axi_conv_knl_RRESP        ( m_axi_RRESP  [2] )
        , .m_axi_conv_knl_RLAST        ( m_axi_RLAST  [2] )
        , .m_axi_conv_knl_RVALID       ( m_axi_RVALID [2] )
        , .m_axi_conv_knl_RREADY       ( m_axi_RREADY [2] )

        , .m_axi_conv_ftu_AWID         ( m_axi_AWID   [3] )
        , .m_axi_conv_ftu_AWADDR       ( m_axi_AWADDR [3] )
        , .m_axi_conv_ftu_AWLEN        ( m_axi_AWLEN  [3] )
        , .m_axi_conv_ftu_AWSIZE       ( m_axi_AWSIZE [3] )
        , .m_axi_conv_ftu_AWBURST      ( m_axi_AWBURST[3] )
        , .m_axi_conv_ftu_AWVALID      ( m_axi_AWVALID[3] )
        , .m_axi_conv_ftu_AWREADY      ( m_axi_AWREADY[3] )
        , .m_axi_conv_ftu_WDATA        ( m_axi_WDATA  [3] )
        , .m_axi_conv_ftu_WSTRB        ( m_axi_WSTRB  [3] )
        , .m_axi_conv_ftu_WLAST        ( m_axi_WLAST  [3] )
        , .m_axi_conv_ftu_WVALID       ( m_axi_WVALID [3] )
        , .m_axi_conv_ftu_WREADY       ( m_axi_WREADY [3] )
        , .m_axi_conv_ftu_BID          ( m_axi_BID    [3] )
        , .m_axi_conv_ftu_BRESP        ( m_axi_BRESP  [3] )
        , .m_axi_conv_ftu_BVALID       ( m_axi_BVALID [3] )
        , .m_axi_conv_ftu_BREADY       ( m_axi_BREADY [3] )
        , .m_axi_conv_ftu_ARID         ( m_axi_ARID   [3] )
        , .m_axi_conv_ftu_ARADDR       ( m_axi_ARADDR [3] )
        , .m_axi_conv_ftu_ARLEN        ( m_axi_ARLEN  [3] )
        , .m_axi_conv_ftu_ARSIZE       ( m_axi_ARSIZE [3] )
        , .m_axi_conv_ftu_ARBURST      ( m_axi_ARBURST[3] )
        , .m_axi_conv_ftu_ARVALID      ( m_axi_ARVALID[3] )
        , .m_axi_conv_ftu_ARREADY      ( m_axi_ARREADY[3] )
        , .m_axi_conv_ftu_RID          ( m_axi_RID    [3] )
        , .m_axi_conv_ftu_RDATA        ( m_axi_RDATA  [3] )
        , .m_axi_conv_ftu_RRESP        ( m_axi_RRESP  [3] )
        , .m_axi_conv_ftu_RLAST        ( m_axi_RLAST  [3] )
        , .m_axi_conv_ftu_RVALID       ( m_axi_RVALID [3] )
        , .m_axi_conv_ftu_RREADY       ( m_axi_RREADY [3] )

        , .interrupt_conv              (  )

        , .m_axi_pool_AWID             ( m_axi_AWID   [4] )
        , .m_axi_pool_AWADDR           ( m_axi_AWADDR [4] )
        , .m_axi_pool_AWLEN            ( m_axi_AWLEN  [4] )
        , .m_axi_pool_AWSIZE           ( m_axi_AWSIZE [4] )
        , .m_axi_pool_AWBURST          ( m_axi_AWBURST[4] )
        , .m_axi_pool_AWVALID          ( m_axi_AWVALID[4] )
        , .m_axi_pool_AWREADY          ( m_axi_AWREADY[4] )
        , .m_axi_pool_WDATA            ( m_axi_WDATA  [4] )
        , .m_axi_pool_WSTRB            ( m_axi_WSTRB  [4] )
        , .m_axi_pool_WLAST            ( m_axi_WLAST  [4] )
        , .m_axi_pool_WVALID           ( m_axi_WVALID [4] )
        , .m_axi_pool_WREADY           ( m_axi_WREADY [4] )
        , .m_axi_pool_BID              ( m_axi_BID    [4] )
        , .m_axi_pool_BRESP            ( m_axi_BRESP  [4] )
        , .m_axi_pool_BVALID           ( m_axi_BVALID [4] )
        , .m_axi_pool_BREADY           ( m_axi_BREADY [4] )
        , .m_axi_pool_ARID             ( m_axi_ARID   [4] )
        , .m_axi_pool_ARADDR           ( m_axi_ARADDR [4] )
        , .m_axi_pool_ARLEN            ( m_axi_ARLEN  [4] )
        , .m_axi_pool_ARSIZE           ( m_axi_ARSIZE [4] )
        , .m_axi_pool_ARBURST          ( m_axi_ARBURST[4] )
        , .m_axi_pool_ARVALID          ( m_axi_ARVALID[4] )
        , .m_axi_pool_ARREADY          ( m_axi_ARREADY[4] )
        , .m_axi_pool_RID              ( m_axi_RID    [4] )
        , .m_axi_pool_RDATA            ( m_axi_RDATA  [4] )
        , .m_axi_pool_RRESP            ( m_axi_RRESP  [4] )
        , .m_axi_pool_RLAST            ( m_axi_RLAST  [4] )
        , .m_axi_pool_RVALID           ( m_axi_RVALID [4] )
        , .m_axi_pool_RREADY           ( m_axi_RREADY [4] )

        , .interrupt_pool              (  )

        , .m_axi_linear_rst_AWID       ( m_axi_AWID   [5] )
        , .m_axi_linear_rst_AWADDR     ( m_axi_AWADDR [5] )
        , .m_axi_linear_rst_AWLEN      ( m_axi_AWLEN  [5] )
        , .m_axi_linear_rst_AWSIZE     ( m_axi_AWSIZE [5] )
        , .m_axi_linear_rst_AWBURST    ( m_axi_AWBURST[5] )
        , .m_axi_linear_rst_AWVALID    ( m_axi_AWVALID[5] )
        , .m_axi_linear_rst_AWREADY    ( m_axi_AWREADY[5] )
        , .m_axi_linear_rst_WDATA      ( m_axi_WDATA  [5] )
        , .m_axi_linear_rst_WSTRB      ( m_axi_WSTRB  [5] )
        , .m_axi_linear_rst_WLAST      ( m_axi_WLAST  [5] )
        , .m_axi_linear_rst_WVALID     ( m_axi_WVALID [5] )
        , .m_axi_linear_rst_WREADY     ( m_axi_WREADY [5] )
        , .m_axi_linear_rst_BID        ( m_axi_BID    [5] )
        , .m_axi_linear_rst_BRESP      ( m_axi_BRESP  [5] )
        , .m_axi_linear_rst_BVALID     ( m_axi_BVALID [5] )
        , .m_axi_linear_rst_BREADY     ( m_axi_BREADY [5] )
        , .m_axi_linear_rst_ARID       ( m_axi_ARID   [5] )
        , .m_axi_linear_rst_ARADDR     ( m_axi_ARADDR [5] )
        , .m_axi_linear_rst_ARLEN      ( m_axi_ARLEN  [5] )
        , .m_axi_linear_rst_ARSIZE     ( m_axi_ARSIZE [5] )
        , .m_axi_linear_rst_ARBURST    ( m_axi_ARBURST[5] )
        , .m_axi_linear_rst_ARVALID    ( m_axi_ARVALID[5] )
        , .m_axi_linear_rst_ARREADY    ( m_axi_ARREADY[5] )
        , .m_axi_linear_rst_RID        ( m_axi_RID    [5] )
        , .m_axi_linear_rst_RDATA      ( m_axi_RDATA  [5] )
        , .m_axi_linear_rst_RRESP      ( m_axi_RRESP  [5] )
        , .m_axi_linear_rst_RLAST      ( m_axi_RLAST  [5] )
        , .m_axi_linear_rst_RVALID     ( m_axi_RVALID [5] )
        , .m_axi_linear_rst_RREADY     ( m_axi_RREADY [5] )

        , .m_axi_linear_weight_AWID    ( m_axi_AWID   [6] )
        , .m_axi_linear_weight_AWADDR  ( m_axi_AWADDR [6] )
        , .m_axi_linear_weight_AWLEN   ( m_axi_AWLEN  [6] )
        , .m_axi_linear_weight_AWSIZE  ( m_axi_AWSIZE [6] )
        , .m_axi_linear_weight_AWBURST ( m_axi_AWBURST[6] )
        , .m_axi_linear_weight_AWVALID ( m_axi_AWVALID[6] )
        , .m_axi_linear_weight_AWREADY ( m_axi_AWREADY[6] )
        , .m_axi_linear_weight_WDATA   ( m_axi_WDATA  [6] )
        , .m_axi_linear_weight_WSTRB   ( m_axi_WSTRB  [6] )
        , .m_axi_linear_weight_WLAST   ( m_axi_WLAST  [6] )
        , .m_axi_linear_weight_WVALID  ( m_axi_WVALID [6] )
        , .m_axi_linear_weight_WREADY  ( m_axi_WREADY [6] )
        , .m_axi_linear_weight_BID     ( m_axi_BID    [6] )
        , .m_axi_linear_weight_BRESP   ( m_axi_BRESP  [6] )
        , .m_axi_linear_weight_BVALID  ( m_axi_BVALID [6] )
        , .m_axi_linear_weight_BREADY  ( m_axi_BREADY [6] )
        , .m_axi_linear_weight_ARID    ( m_axi_ARID   [6] )
        , .m_axi_linear_weight_ARADDR  ( m_axi_ARADDR [6] )
        , .m_axi_linear_weight_ARLEN   ( m_axi_ARLEN  [6] )
        , .m_axi_linear_weight_ARSIZE  ( m_axi_ARSIZE [6] )
        , .m_axi_linear_weight_ARBURST ( m_axi_ARBURST[6] )
        , .m_axi_linear_weight_ARVALID ( m_axi_ARVALID[6] )
        , .m_axi_linear_weight_ARREADY ( m_axi_ARREADY[6] )
        , .m_axi_linear_weight_RID     ( m_axi_RID    [6] )
        , .m_axi_linear_weight_RDATA   ( m_axi_RDATA  [6] )
        , .m_axi_linear_weight_RRESP   ( m_axi_RRESP  [6] )
        , .m_axi_linear_weight_RLAST   ( m_axi_RLAST  [6] )
        , .m_axi_linear_weight_RVALID  ( m_axi_RVALID [6] )
        , .m_axi_linear_weight_RREADY  ( m_axi_RREADY [6] )

        , .interrupt_linear            (  )

        , .m_axi_mover_AWID            ( m_axi_AWID   [7] )
        , .m_axi_mover_AWADDR          ( m_axi_AWADDR [7] )
        , .m_axi_mover_AWLEN           ( m_axi_AWLEN  [7] )
        , .m_axi_mover_AWSIZE          ( m_axi_AWSIZE [7] )
        , .m_axi_mover_AWBURST         ( m_axi_AWBURST[7] )
        , .m_axi_mover_AWVALID         ( m_axi_AWVALID[7] )
        , .m_axi_mover_AWREADY         ( m_axi_AWREADY[7] )
        , .m_axi_mover_WDATA           ( m_axi_WDATA  [7] )
        , .m_axi_mover_WSTRB           ( m_axi_WSTRB  [7] )
        , .m_axi_mover_WLAST           ( m_axi_WLAST  [7] )
        , .m_axi_mover_WVALID          ( m_axi_WVALID [7] )
        , .m_axi_mover_WREADY          ( m_axi_WREADY [7] )
        , .m_axi_mover_BID             ( m_axi_BID    [7] )
        , .m_axi_mover_BRESP           ( m_axi_BRESP  [7] )
        , .m_axi_mover_BVALID          ( m_axi_BVALID [7] )
        , .m_axi_mover_BREADY          ( m_axi_BREADY [7] )
        , .m_axi_mover_ARID            ( m_axi_ARID   [7] )
        , .m_axi_mover_ARADDR          ( m_axi_ARADDR [7] )
        , .m_axi_mover_ARLEN           ( m_axi_ARLEN  [7] )
        , .m_axi_mover_ARSIZE          ( m_axi_ARSIZE [7] )
        , .m_axi_mover_ARBURST         ( m_axi_ARBURST[7] )
        , .m_axi_mover_ARVALID         ( m_axi_ARVALID[7] )
        , .m_axi_mover_ARREADY         ( m_axi_ARREADY[7] )
        , .m_axi_mover_RID             ( m_axi_RID    [7] )
        , .m_axi_mover_RDATA           ( m_axi_RDATA  [7] )
        , .m_axi_mover_RRESP           ( m_axi_RRESP  [7] )
        , .m_axi_mover_RLAST           ( m_axi_RLAST  [7] )
        , .m_axi_mover_RVALID          ( m_axi_RVALID [7] )
        , .m_axi_mover_RREADY          ( m_axi_RREADY [7] )

        , .interrupt_mover             (  )
    );

    assign m_axi_ARLOCK={P_NUM_AXI_MASTER{1'b0}};
    assign m_axi_AWLOCK={P_NUM_AXI_MASTER{1'b0}};
